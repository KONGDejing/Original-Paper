`timescale 1ns/1ps
module sram_test_fangxin
(
    input CLK,     //120M
	 input RSTn,
	 
	 input PCLK,
	 input HREF,
	 input VSYNC_ov7620_L,
	 input [7:0]Y_Data,

	 output[17:0]sram_addr,
	 output sram_wr_n,
	 output sram_ce_n,
	 inout[7:0]sram_data,
	 
	 output HSYNC,
    output VSYNC,
	 output [2:0]RGB_Sig
);

/*******************VGAͬ��****************************/

reg [10:0]C1;
reg [9:0]C2;
reg rH,rV;
reg sram_ce_r; 
	 always @ ( posedge CLK or negedge RSTn )
	     if( !RSTn )
		      begin
				    C1 <= 11'd0;
					 C2 <= 10'd0;
					 rH <= 1'b1;
					 rV <= 1'b1;
					 sram_ce_r<=1'b1;
				end
		  else 
		      begin
				    
					 if( C1 == 1904 ) rH <= 1'b0; 
				     else if( C1 == 152  ) rH <= 1'b1;
				     //else if( C1 == 0 ) rH <= 1'b0;
					 
					 if( C2 == 932 ) rV <= 1'b0;
					 else if( C2 == 3  ) rV <= 1'b1;
					 //else if( C2 == 0 ) rV <= 1'b0;
					 
					 if( C2 == 932 ) C2 <= 10'd1;
					 else if( C1 == 1904 ) C2 <= C2 + 1'b1;
					 
				     if( C1 == 1904 ) C1 <= 11'd1;
					 else C1 <= C1 + 1'b1;
					 
					 sram_ce_r<=1'b0;
					 
				end
assign HSYNC = rH;
assign VSYNC = rV;
assign sram_ce_n=sram_ce_r;	 
//-----------------------------------------------------------
/********************VGAɨ��*********************************/
	 
	 parameter _X = 10'd640, _Y = 10'd240, _XOFF = 10'd0, _YOFF = 10'd25; 
	 
/**************************************/
    reg isRectangle;
    reg [17:0]x,y;
	 reg [17:0]ADDR_R;


    always @ ( posedge CLK or negedge RSTn )
	     if( !RSTn )
		      begin
				    x <= 18'd0;
					 y <= 18'd0;
				    ADDR_R<=18'd0;
				  
				end
			else
			   begin
				
				    // step 1 : compute data address and index-n
					 if( (C1 > 152 + 232 + _XOFF && C1 <= 152 + 232 + _XOFF +_X) && 
					     (C2 > 3 + 28 + _YOFF && C2 <= 3 + 28 + _YOFF + _Y) && VGA_r)
					     begin 
						      isRectangle <= 1'b1;
						      x <= C1 - _XOFF - 152 - 232 - 1; 
						      y <= C2 - _YOFF - 3 - 28 - 1;
					         ADDR_R = (y << 9 +  y <<7) + x ; //address = y*640+x
					     end
						 
					 else 
					         isRectangle <= 1'b0;
		       end
/*****************************************************/

reg [7:0]wr_data;
reg [7:0]rd_data;
reg [17:0]addr_r;
reg [3:0]i;

wire sram_wr_req;
wire sram_rd_req;
reg VGA_r,Collect_r;
always @(posedge CLK or negedge RSTn)
     if(!RSTn)
		   begin
				 i<=4'd0;  
				 VGA_r<=1'd0;
				 Collect_r<=1'd0;
			end
		 else 
		   case(i)
			   0:
				if(VSYNC_ov7620_L)begin  i<=1'b1;   end
				else
			   	begin
						  VGA_r<=1'd0;
						  Collect_r<=1'd1; 
				   end
	         1,2,3:
		   	if(VSYNC_ov7620_L)begin  i<=i+1'b1; end
				else
					begin
					     VGA_r<=1'd1;
						  Collect_r<=1'd0;
					end
				4:      begin  i<=4'd0;  end 
			 endcase
//---------------------------------------------------
reg sram_wr_req_r;
reg [1:0]j;
always @(posedge PCLK or negedge RSTn)           //or negedge RSTn and Collect_r
   if(!RSTn)sram_wr_req_r<=1'b0;
   else
	begin
		 if(~VSYNC_ov7620_L)
			 begin 
				 if(HREF & Collect_r)
				      begin
								 case(j)
									 0:begin sram_wr_req_r<=1'b1;j<=j+1'b1; end
									 1:begin sram_wr_req_r<=1'b0;j<=1'b0; end
								 endcase
						end		
				 else
				     sram_wr_req_r<=1'b0;
			 end
		 else
		    sram_wr_req_r<=1'b0;
	end  
assign sram_wr_req=sram_wr_req_r;
assign sram_rd_req=(ADDR_R%2==1);

always @(posedge CLK or negedge RSTn)
     if(!RSTn)begin addr_r<=18'd0;end	    
	  else if(sram_wr_req) begin addr_r<=addr_r+1'b1; end
	  
assign sram_addr=Collect_r ? addr_r : ADDR_R;

//-------------------------------------------------

`define DELAY_20NS    (cnt==3'd1)
reg [2:0]cnt;

always @(posedge CLK or negedge RSTn)
     if(!RSTn) cnt<=3'd0;
     else if(cstate==IDLE)cnt<=3'd0;
	  else cnt<=cnt+1'b1;
	  
//------------------����ʽ״̬��-------------------------------
parameter IDLE =4'd0,
          WRT0 =4'd1,
			 WRT1 =4'd2,
			 REA0 =4'd3,
			 REA1 =4'd4;
reg [3:0]cstate,nstate;

always @(posedge CLK or negedge RSTn)
    if(!RSTn)cstate<=IDLE;
	 else cstate<=nstate;
	 
always @(cstate or sram_wr_req or sram_rd_req or cnt)
    case(cstate)
	      IDLE: if(sram_wr_req)nstate<=WRT0;
			      else if(sram_rd_req)nstate<=REA0;
					else nstate<=IDLE;
			WRT0: if(`DELAY_20NS) nstate<=WRT1;
			      else nstate<=WRT0;
			WRT1: nstate<=IDLE;
			REA0: if(`DELAY_20NS) nstate<=REA1;
			      else nstate<=REA0;
			REA1: nstate<=IDLE;
		default: nstate<=IDLE;
	endcase
			 
//------------------------------------------------
//always @(posedge CLK or negedge RSTn)
//    if(!RSTn)wr_data<=8'd0;
//	 else if(cstate==WRT1)wr_data<=Y_Data;

reg sdlink;
	
always @(posedge CLK or negedge RSTn)
    if(!RSTn)sdlink<=1'b0;
	 else
	    case(cstate)
		     IDLE: if(sram_wr_req)sdlink <=1'b1;
			        else if(sram_rd_req)sdlink<=1'b0;
					  else sdlink<=1'b0;
			  WRT0: sdlink<=1'b1;
			  default: sdlink<=1'b0;
			  endcase
			  
assign sram_data = sdlink ? Y_Data : 8'hzz;       //д����
assign sram_wr_n = ~sdlink;

always @(posedge CLK or negedge RSTn)
    if(!RSTn)rd_data<=8'd0;
    else if(cstate==REA1)rd_data<=sram_data;	     //������
//---------------------------------------------------	 
reg [2:0]rRGB;
always @ (posedge CLK or negedge RSTn)
         if(!RSTn)
			       rRGB<=3'b000;
         else if(VGA_r)
						begin			
							   if(rd_data<=8'b01111110)
										 rRGB<=3'b000;
								else			 
										 rRGB<=3'b111;
						end
			else
			 rRGB<=3'b000; 
			
/*******************************************************/

assign RGB_Sig=( isRectangle && VGA_r)? rRGB : 3'b000;
		  
endmodule


